--library IEEE;
--use IEEE.std_logic_1164.all;

entity temp is
  port (A: in bit;
        Y: out bit);
end temp;

architecture behave of temp is
constant c : bit := '1';
begin
  y <= a;

end behave;        
